`timescale 1ns/1ps

module Controller();
    //
endmodule
